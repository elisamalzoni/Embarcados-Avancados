-- unsaved_tb.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity unsaved_tb is
end entity unsaved_tb;

architecture rtl of unsaved_tb is
	component unsaved is
		port (
			clk_clk                   : in  std_logic                    := 'X';             -- clk
			key_export                : in  std_logic_vector(3 downto 0) := (others => 'X'); -- export
			leds_writeresponsevalid_n : out std_logic_vector(3 downto 0);                    -- writeresponsevalid_n
			reset_reset_n             : in  std_logic                    := 'X'              -- reset_n
		);
	end component unsaved;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_conduit_bfm is
		port (
			sig_export : out std_logic_vector(3 downto 0)   -- export
		);
	end component altera_conduit_bfm;

	component altera_conduit_bfm_0002 is
		port (
			clk                      : in std_logic                    := 'X';             -- clk
			sig_writeresponsevalid_n : in std_logic_vector(3 downto 0) := (others => 'X'); -- writeresponsevalid_n
			reset                    : in std_logic                    := 'X'              -- reset
		);
	end component altera_conduit_bfm_0002;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal unsaved_inst_clk_bfm_clk_clk           : std_logic;                    -- unsaved_inst_clk_bfm:clk -> [unsaved_inst:clk_clk, unsaved_inst_leds_bfm:clk, unsaved_inst_reset_bfm:clk]
	signal unsaved_inst_key_bfm_conduit_export    : std_logic_vector(3 downto 0); -- unsaved_inst_key_bfm:sig_export -> unsaved_inst:key_export
	signal unsaved_inst_leds_writeresponsevalid_n : std_logic_vector(3 downto 0); -- unsaved_inst:leds_writeresponsevalid_n -> unsaved_inst_leds_bfm:sig_writeresponsevalid_n
	signal unsaved_inst_reset_bfm_reset_reset     : std_logic;                    -- unsaved_inst_reset_bfm:reset -> unsaved_inst:reset_reset_n

begin

	unsaved_inst : component unsaved
		port map (
			clk_clk                   => unsaved_inst_clk_bfm_clk_clk,           --   clk.clk
			key_export                => unsaved_inst_key_bfm_conduit_export,    --   key.export
			leds_writeresponsevalid_n => unsaved_inst_leds_writeresponsevalid_n, --  leds.writeresponsevalid_n
			reset_reset_n             => unsaved_inst_reset_bfm_reset_reset      -- reset.reset_n
		);

	unsaved_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => unsaved_inst_clk_bfm_clk_clk  -- clk.clk
		);

	unsaved_inst_key_bfm : component altera_conduit_bfm
		port map (
			sig_export => unsaved_inst_key_bfm_conduit_export  -- conduit.export
		);

	unsaved_inst_leds_bfm : component altera_conduit_bfm_0002
		port map (
			clk                      => unsaved_inst_clk_bfm_clk_clk,           --     clk.clk
			sig_writeresponsevalid_n => unsaved_inst_leds_writeresponsevalid_n, -- conduit.writeresponsevalid_n
			reset                    => '0'                                     -- (terminated)
		);

	unsaved_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => unsaved_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => unsaved_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of unsaved_tb
